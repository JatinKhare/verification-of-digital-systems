module seq_top ( );
    mul  spec( );
    mul  impl( );
endmodule

