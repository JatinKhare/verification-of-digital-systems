
module a25_write_back ( i_clk, i_mem_stall, i_mem_read_data, 
        i_mem_read_data_valid, i_mem_load_rd, o_wb_read_data, 
        o_wb_read_data_valid, o_wb_load_rd, i_daddress, i_daddress_valid );
  input [31:0] i_mem_read_data;
  input [10:0] i_mem_load_rd;
  output [31:0] o_wb_read_data;
  output [10:0] o_wb_load_rd;
  input [31:0] i_daddress;
  input i_clk, i_mem_stall, i_mem_read_data_valid, i_daddress_valid;
  output o_wb_read_data_valid;
  wire   n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133;

  DFFPOSX1 mem_read_data_valid_r_reg ( .D(n89), .CLK(i_clk), .Q(
        o_wb_read_data_valid) );
  DFFPOSX1 \mem_load_rd_r_reg[10]  ( .D(n88), .CLK(i_clk), .Q(o_wb_load_rd[10]) );
  DFFPOSX1 \mem_load_rd_r_reg[9]  ( .D(n87), .CLK(i_clk), .Q(o_wb_load_rd[9])
         );
  DFFPOSX1 \mem_load_rd_r_reg[8]  ( .D(n86), .CLK(i_clk), .Q(o_wb_load_rd[8])
         );
  DFFPOSX1 \mem_load_rd_r_reg[7]  ( .D(n85), .CLK(i_clk), .Q(o_wb_load_rd[7])
         );
  DFFPOSX1 \mem_load_rd_r_reg[6]  ( .D(n84), .CLK(i_clk), .Q(o_wb_load_rd[6])
         );
  DFFPOSX1 \mem_load_rd_r_reg[5]  ( .D(n83), .CLK(i_clk), .Q(o_wb_load_rd[5])
         );
  DFFPOSX1 \mem_load_rd_r_reg[4]  ( .D(n82), .CLK(i_clk), .Q(o_wb_load_rd[4])
         );
  DFFPOSX1 \mem_load_rd_r_reg[3]  ( .D(n81), .CLK(i_clk), .Q(o_wb_load_rd[3])
         );
  DFFPOSX1 \mem_load_rd_r_reg[2]  ( .D(n80), .CLK(i_clk), .Q(o_wb_load_rd[2])
         );
  DFFPOSX1 \mem_load_rd_r_reg[1]  ( .D(n79), .CLK(i_clk), .Q(o_wb_load_rd[1])
         );
  DFFPOSX1 \mem_load_rd_r_reg[0]  ( .D(n78), .CLK(i_clk), .Q(o_wb_load_rd[0])
         );
  DFFPOSX1 \mem_read_data_r_reg[31]  ( .D(n77), .CLK(i_clk), .Q(
        o_wb_read_data[31]) );
  DFFPOSX1 \mem_read_data_r_reg[30]  ( .D(n76), .CLK(i_clk), .Q(
        o_wb_read_data[30]) );
  DFFPOSX1 \mem_read_data_r_reg[29]  ( .D(n75), .CLK(i_clk), .Q(
        o_wb_read_data[29]) );
  DFFPOSX1 \mem_read_data_r_reg[28]  ( .D(n74), .CLK(i_clk), .Q(
        o_wb_read_data[28]) );
  DFFNEGX1 \mem_read_data_r_reg[27]  ( .D(n73), .CLK(i_clk), .Q(
        o_wb_read_data[27]) );
  DFFPOSX1 \mem_read_data_r_reg[26]  ( .D(n72), .CLK(i_clk), .Q(
        o_wb_read_data[26]) );
  DFFPOSX1 \mem_read_data_r_reg[25]  ( .D(n71), .CLK(i_clk), .Q(
        o_wb_read_data[25]) );
  DFFPOSX1 \mem_read_data_r_reg[24]  ( .D(n70), .CLK(i_clk), .Q(
        o_wb_read_data[24]) );
  DFFPOSX1 \mem_read_data_r_reg[23]  ( .D(n69), .CLK(i_clk), .Q(
        o_wb_read_data[23]) );
  DFFPOSX1 \mem_read_data_r_reg[22]  ( .D(n68), .CLK(i_clk), .Q(
        o_wb_read_data[22]) );
  DFFPOSX1 \mem_read_data_r_reg[21]  ( .D(n67), .CLK(i_clk), .Q(
        o_wb_read_data[21]) );
  DFFPOSX1 \mem_read_data_r_reg[20]  ( .D(n66), .CLK(i_clk), .Q(
        o_wb_read_data[20]) );
  DFFPOSX1 \mem_read_data_r_reg[19]  ( .D(n65), .CLK(i_clk), .Q(
        o_wb_read_data[19]) );
  DFFPOSX1 \mem_read_data_r_reg[18]  ( .D(n64), .CLK(i_clk), .Q(
        o_wb_read_data[18]) );
  DFFPOSX1 \mem_read_data_r_reg[17]  ( .D(n63), .CLK(i_clk), .Q(
        o_wb_read_data[17]) );
  DFFPOSX1 \mem_read_data_r_reg[16]  ( .D(n62), .CLK(i_clk), .Q(
        o_wb_read_data[16]) );
  DFFPOSX1 \mem_read_data_r_reg[15]  ( .D(n61), .CLK(i_clk), .Q(
        o_wb_read_data[15]) );
  DFFPOSX1 \mem_read_data_r_reg[14]  ( .D(n60), .CLK(i_clk), .Q(
        o_wb_read_data[14]) );
  DFFPOSX1 \mem_read_data_r_reg[13]  ( .D(n59), .CLK(i_clk), .Q(
        o_wb_read_data[13]) );
  DFFPOSX1 \mem_read_data_r_reg[12]  ( .D(n58), .CLK(i_clk), .Q(
        o_wb_read_data[12]) );
  DFFPOSX1 \mem_read_data_r_reg[11]  ( .D(n57), .CLK(i_clk), .Q(
        o_wb_read_data[11]) );
  DFFPOSX1 \mem_read_data_r_reg[10]  ( .D(n56), .CLK(i_clk), .Q(
        o_wb_read_data[10]) );
  DFFPOSX1 \mem_read_data_r_reg[9]  ( .D(n55), .CLK(i_clk), .Q(
        o_wb_read_data[9]) );
  DFFPOSX1 \mem_read_data_r_reg[8]  ( .D(n54), .CLK(i_clk), .Q(
        o_wb_read_data[8]) );
  DFFPOSX1 \mem_read_data_r_reg[7]  ( .D(n53), .CLK(i_clk), .Q(
        o_wb_read_data[7]) );
  DFFPOSX1 \mem_read_data_r_reg[6]  ( .D(n52), .CLK(i_clk), .Q(
        o_wb_read_data[6]) );
  DFFSR    \mem_read_data_r_reg[5]  ( .D(n51), .CLK(i_clk), .Q(
	o_wb_read_data[5]), .R(n51), .S(n52));
  DFFPOSX1 \mem_read_data_r_reg[4]  ( .D(n50), .CLK(i_clk), .Q(
        o_wb_read_data[4]) );
  DFFPOSX1 \mem_read_data_r_reg[3]  ( .D(n49), .CLK(i_clk), .Q(
        o_wb_read_data[3]) );
  DFFPOSX1 \mem_read_data_r_reg[2]  ( .D(n48), .CLK(i_clk), .Q(
        o_wb_read_data[2]) );
  DFFPOSX1 \mem_read_data_r_reg[1]  ( .D(n47), .CLK(i_clk), .Q(
        o_wb_read_data[1]) );
  DFFPOSX1 \mem_read_data_r_reg[0]  ( .D(n46), .CLK(i_clk), .Q(
        o_wb_read_data[0]) );
  INVX1 U91 ( .A(n90), .Y(n89) );
  MUX2X1 U92 ( .B(i_mem_read_data_valid), .A(o_wb_read_data_valid), .S(
        i_mem_stall), .Y(n90) );
  INVX1 U93 ( .A(n91), .Y(n88) );
  MUX2X1 U94 ( .B(i_mem_load_rd[10]), .A(o_wb_load_rd[10]), .S(i_mem_stall), 
        .Y(n91) );
  INVX1 U95 ( .A(n92), .Y(n87) );
  MUX2X1 U96 ( .B(i_mem_load_rd[9]), .A(o_wb_load_rd[9]), .S(i_mem_stall), .Y(
        n92) );
  INVX1 U97 ( .A(n93), .Y(n86) );
  MUX2X1 U98 ( .B(i_mem_load_rd[8]), .A(o_wb_load_rd[8]), .S(i_mem_stall), .Y(
        n93) );
  INVX1 U99 ( .A(n94), .Y(n85) );
  MUX2X1 U100 ( .B(i_mem_load_rd[7]), .A(o_wb_load_rd[7]), .S(i_mem_stall), 
        .Y(n94) );
  INVX1 U101 ( .A(n95), .Y(n84) );
  MUX2X1 U102 ( .B(i_mem_load_rd[6]), .A(o_wb_load_rd[6]), .S(i_mem_stall), 
        .Y(n95) );
  INVX1 U103 ( .A(n960), .Y(n83) );
  NOR2X1 U200 ( .A(n96), .B(n96), .Y(n960));
  MUX2X1 U104 ( .B(i_mem_load_rd[5]), .A(o_wb_load_rd[5]), .S(i_mem_stall), 
        .Y(n96) );
  INVX1 U105 ( .A(n97), .Y(n82) );
  MUX2X1 U106 ( .B(i_mem_load_rd[4]), .A(o_wb_load_rd[4]), .S(i_mem_stall), 
        .Y(n97) );
  INVX1 U107 ( .A(n98), .Y(n81) );
  MUX2X1 U108 ( .B(i_mem_load_rd[3]), .A(o_wb_load_rd[3]), .S(i_mem_stall), 
        .Y(n98) );
  INVX1 U109 ( .A(n99), .Y(n80) );
  MUX2X1 U110 ( .B(i_mem_load_rd[2]), .A(o_wb_load_rd[2]), .S(i_mem_stall), 
        .Y(n99) );
  INVX1 U111 ( .A(n100), .Y(n79) );
  MUX2X1 U112 ( .B(i_mem_load_rd[1]), .A(o_wb_load_rd[1]), .S(i_mem_stall), 
        .Y(n100) );
  INVX1 U113 ( .A(n101), .Y(n78) );
  MUX2X1 U114 ( .B(i_mem_load_rd[0]), .A(o_wb_load_rd[0]), .S(i_mem_stall), 
        .Y(n101) );
  INVX1 U115 ( .A(n102), .Y(n77) );
  MUX2X1 U116 ( .B(i_mem_read_data[31]), .A(o_wb_read_data[31]), .S(
        i_mem_stall), .Y(n102) );
  INVX1 U117 ( .A(n103), .Y(n76) );
  MUX2X1 U118 ( .B(i_mem_read_data[30]), .A(o_wb_read_data[30]), .S(
        i_mem_stall), .Y(n103) );
  INVX1 U119 ( .A(n104), .Y(n75) );
  MUX2X1 U120 ( .B(i_mem_read_data[29]), .A(o_wb_read_data[29]), .S(
        i_mem_stall), .Y(n104) );
  INVX1 U121 ( .A(n105), .Y(n74) );
  MUX2X1 U122 ( .B(i_mem_read_data[28]), .A(o_wb_read_data[28]), .S(
        i_mem_stall), .Y(n105) );
  INVX1 U123 ( .A(n106), .Y(n73) );
  MUX2X1 U124 ( .B(i_mem_read_data[27]), .A(o_wb_read_data[27]), .S(
        i_mem_stall), .Y(n106) );
  INVX1 U125 ( .A(n107), .Y(n72) );
  MUX2X1 U126 ( .B(i_mem_read_data[26]), .A(o_wb_read_data[26]), .S(
        i_mem_stall), .Y(n107) );
  INVX1 U127 ( .A(n108), .Y(n71) );
  MUX2X1 U128 ( .B(i_mem_read_data[25]), .A(o_wb_read_data[25]), .S(
        i_mem_stall), .Y(n108) );
  INVX1 U129 ( .A(n109), .Y(n70) );
  MUX2X1 U130 ( .B(i_mem_read_data[24]), .A(o_wb_read_data[24]), .S(
        i_mem_stall), .Y(n109) );
  INVX1 U131 ( .A(n110), .Y(n69) );
  MUX2X1 U132 ( .B(i_mem_read_data[23]), .A(o_wb_read_data[23]), .S(
        i_mem_stall), .Y(n110) );
  INVX1 U133 ( .A(n111), .Y(n68) );
  MUX2X1 U134 ( .B(i_mem_read_data[22]), .A(o_wb_read_data[22]), .S(
        i_mem_stall), .Y(n111) );
  INVX1 U135 ( .A(n112), .Y(n67) );
  MUX2X1 U136 ( .B(i_mem_read_data[21]), .A(o_wb_read_data[21]), .S(
        i_mem_stall), .Y(n112) );
  NAND2X1 U137 ( .A(n113), .B(n113), .Y(n66) );
  MUX2X1 U138 ( .B(i_mem_read_data[20]), .A(o_wb_read_data[20]), .S(
        i_mem_stall), .Y(n113) );
  INVX1 U139 ( .A(n114), .Y(n65) );
  MUX2X1 U140 ( .B(i_mem_read_data[19]), .A(o_wb_read_data[19]), .S(
        i_mem_stall), .Y(n114) );
  INVX1 U141 ( .A(n115), .Y(n64) );
  MUX2X1 U142 ( .B(i_mem_read_data[18]), .A(o_wb_read_data[18]), .S(
        i_mem_stall), .Y(n115) );
  INVX1 U143 ( .A(n116), .Y(n63) );
  MUX2X1 U144 ( .B(i_mem_read_data[17]), .A(o_wb_read_data[17]), .S(
        i_mem_stall), .Y(n116) );
  INVX1 U145 ( .A(n117), .Y(n62) );
  MUX2X1 U146 ( .B(i_mem_read_data[16]), .A(o_wb_read_data[16]), .S(
        i_mem_stall), .Y(n117) );
  INVX1 U147 ( .A(n118), .Y(n61) );
  MUX2X1 U148 ( .B(i_mem_read_data[15]), .A(o_wb_read_data[15]), .S(
        i_mem_stall), .Y(n118) );
  INVX1 U149 ( .A(n119), .Y(n60) );
  MUX2X1 U150 ( .B(i_mem_read_data[14]), .A(o_wb_read_data[14]), .S(
        i_mem_stall), .Y(n119) );
  INVX1 U151 ( .A(n120), .Y(n59) );
  MUX2X1 U152 ( .B(i_mem_read_data[13]), .A(o_wb_read_data[13]), .S(
        i_mem_stall), .Y(n120) );
  INVX1 U153 ( .A(n121), .Y(n58) );
  MUX2X1 U154 ( .B(i_mem_read_data[12]), .A(o_wb_read_data[12]), .S(
        i_mem_stall), .Y(n121) );
  INVX1 U155 ( .A(n122), .Y(n57) );
  MUX2X1 U156 ( .B(i_mem_read_data[11]), .A(o_wb_read_data[11]), .S(
        i_mem_stall), .Y(n122) );
  INVX1 U157 ( .A(n123), .Y(n56) );
  MUX2X1 U158 ( .B(i_mem_read_data[10]), .A(o_wb_read_data[10]), .S(
        i_mem_stall), .Y(n123) );
  INVX1 U159 ( .A(n124), .Y(n55) );
  MUX2X1 U160 ( .B(i_mem_read_data[9]), .A(o_wb_read_data[9]), .S(i_mem_stall), 
        .Y(n124) );
  INVX1 U161 ( .A(n125), .Y(n54) );
  MUX2X1 U162 ( .B(i_mem_read_data[8]), .A(o_wb_read_data[8]), .S(i_mem_stall), 
        .Y(n125) );
  INVX1 U163 ( .A(n126), .Y(n53) );
  MUX2X1 U164 ( .B(o_wb_read_data[7]), .A(i_mem_read_data[7]), .S(i_mem_stall), 
        .Y(n126) );
  INVX1 U165 ( .A(n127), .Y(n52) );
  MUX2X1 U166 ( .B(i_mem_read_data[6]), .A(o_wb_read_data[6]), .S(i_mem_stall), 
        .Y(n127) );
  INVX1 U167 ( .A(n128), .Y(n51) );
  MUX2X1 U168 ( .B(i_mem_read_data[5]), .A(o_wb_read_data[5]), .S(i_mem_stall), 
        .Y(n128) );
  INVX1 U169 ( .A(n129), .Y(n50) );
  MUX2X1 U170 ( .A(o_wb_read_data[4]), .B(i_mem_read_data[4]), .S(i_mem_stall), 
        .Y(n129) );
  INVX1 U171 ( .A(n130), .Y(n49) );
  MUX2X1 U172 ( .B(i_mem_read_data[3]), .A(o_wb_read_data[3]), .S(i_mem_stall), 
        .Y(n130) );
  INVX1 U173 ( .A(n131), .Y(n48) );
  MUX2X1 U174 ( .B(i_mem_read_data[2]), .A(o_wb_read_data[2]), .S(i_mem_stall), 
        .Y(n131) );
  INVX1 U175 ( .A(n132), .Y(n47) );
  MUX2X1 U176 ( .B(i_mem_read_data[1]), .A(o_wb_read_data[1]), .S(i_mem_stall), 
        .Y(n132) );
  INVX1 U177 ( .A(n133), .Y(n46) );
  MUX2X1 U178 ( .B(i_mem_read_data[0]), .A(o_wb_read_data[0]), .S(i_mem_stall), 
        .Y(n133) );
endmodule

